* MOC3040 TRIAC Circuit Simulation

* Power Supply
V1 1 0 AC 220 50          ; AC mains voltage

* MOC3040 LED Input
R1 2 3 330                ; Current limiting resistor
D1 3 0 LED                ; LED model
V2 2 0 PULSE(0 5 0 1u 1u 10m 20m) ; Input trigger signal

* MOC3040 Phototransistor
Q1 5 4 0 NPN
R2 4 5 1k
V3 4 0 5

* TRIAC Subcircuit Definition
.SUBCKT TRIACMODEL A G K
S1 A G K M1             ; Switch for one polarity
S2 K G A M1             ; Switch for opposite polarity
.MODEL M1 SW (RON=1 ROFF=1MEG VT=1.2 VH=0.1) ; Switch model
.ENDS TRIACMODEL

* TRIAC and Load
XTRIAC 5 6 0 TRIACMODEL   ; TRIAC controlled by MOC3040
R3 6 0 10                 ; Load resistor

* LED Model
.MODEL LED D (IS=1e-14 N=1.5)

* NPN Transistor Model
.MODEL NPN NPN (IS=1e-14 BF=100)

* Simulation Control
.TRAN 0 100m 0 1m
.PLOT TRAN V(6)
.END